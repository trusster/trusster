`include "/users/mmintz/book_install/truss/inc/truss_verification_component.svh"

program killme;

endprogram