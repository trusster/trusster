/*
Trusster Open Source License version 1.0a (TRUST)
copyright (c) 2006 Mike Mintz and Robert Ekendahl.  All rights reserved. 

Redistribution and use in source and binary forms, with or without modification, 
are permitted provided that the following conditions are met: 
   
  * Redistributions of source code must retain the above copyright notice, 
    this list of conditions and the following disclaimer.
  * Redistributions in binary form must reproduce the above copyright notice, 
    this list of conditions and the following disclaimer in the documentation 
    and/or other materials provided with the distribution.
  * Redistributions in any form must be accompanied by information on how to obtain 
    complete source code for this software and any accompanying software that uses this software.
    The source code must either be included in the distribution or be available in a timely fashion for no more than 
    the cost of distribution plus a nominal fee, and must be freely redistributable under reasonable and no more 
    restrictive conditions. For an executable file, complete source code means the source code for all modules it 
    contains. It does not include source code for modules or files that typically accompany the major components 
    of the operating system on which the executable file runs.
 

THIS SOFTWARE IS PROVIDED BY MIKE MINTZ AND ROBERT EKENDAHL ``AS IS'' AND ANY EXPRESS OR IMPLIED WARRANTIES, 
INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE, 
OR NON-INFRINGEMENT, ARE DISCLAIMED. IN NO EVENT SHALL MIKE MINTZ AND ROBERT EKENDAHL OR ITS CONTRIBUTORS 
BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, 
BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; 
OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, 
OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, 
EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
*/
`ifndef __quad_uart_irritators__
`define __quad_uart_irritators__

`include "truss.svh"
`include "testbench.svh"

`include "truss.svh"


  typedef class uart_basic_test_component;
  typedef class uart_basic_irritator;

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
class quad_uart_irritators extends truss::test_base;
   extern function new (testbench tb, truss::watchdog w, string n); 

  extern virtual task time_zero_setup ();
  extern virtual task out_of_reset (truss::reset r);
  extern virtual function void randomize2 ();
  extern virtual task write_to_hardware ();
  extern virtual task start ();
  extern virtual task wait_for_completion ();
  extern virtual function void report (string prefix);
  
  local testbench testbench_;
  local uart_basic_test_component uart_test_component_ingress_;
  local uart_basic_test_component uart_test_component_egress_;

  local uart_basic_irritator uart_basic_irritator_ingress_[number_of_uarts];
  local uart_basic_irritator uart_basic_irritator_egress_[number_of_uarts];


  extern local function void standard_configuration (string name);
  extern local function void standard_generator (string name);

  local rand teal::uint32 uart_index;
  local teal::uint32 min_uart_index;
  local teal::uint32 max_uart_index;
  constraint uart_index_valid {uart_index >= min_uart_index; uart_index <= max_uart_index;}
endclass

`endif
