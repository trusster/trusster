/*
 * Copyright (c) 2004 Mike Mintz (mike@applevalleysoftware.com)
 *
 *    This source code is free software; you can redistribute it
 *    and/or modify it in source code form under the terms of the GNU
 *    General Public License as published by the Free Software
 *    Foundation; either version 2 of the License, or (at your option)
 *    any later version.
 *
 *    This program is distributed in the hope that it will be useful,
 *    but WITHOUT ANY WARRANTY; without even the implied warranty of
 *    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 *    GNU General Public License for more details.
 *
 *    You should have received a copy of the GNU General Public License
 *    along with this program; if not, write to the Free Software
 *    Foundation, Inc., 59 Temple Place - Suite 330, Boston, MA 02111-1307, USA
 */

`timescale 1 ps / 1 ps

module top;
   initial begin
	#10;
	$verification_top;
end

  reg[7:0] run_test;
  initial begin
	run_test = 0;
	#44;
	run_test = 'b1000_0000;
   end

 reg clk;
  initial begin
	clk <= 0;
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
	 #10;
 	  clk <= ~clk; 
$display ("yaya");
  end


endmodule 

