function dictionary_impl::new ();
   //ARRGH because of no statics dictionary cannot have a logger!
   //This is to allow the logger to use the dictionary to see what level the user wants to debug at
   //This log feature is far more important than logger in the dictionary implementtaion class
//   log_ = new ("Dictionary");

endfunction // dictionary_impl

function string dictionary_impl::teal_scan_plusargs (string name);
   string returned;
   bit found = $value$plusargs ({name, "+%s"},returned);
//   $display ("plus args search for %s found %s", name, returned);

  if (found) return returned; else return "";
endfunction 


function string dictionary_impl::find_on_command_line ( string name,  string default_name);
  string arg = teal_scan_plusargs (name);
  return (arg != "") ? arg : default_name;
endfunction



task dictionary_impl::process_file_ (string path);
    integer file_id = $fopen (path, "r");
//   log_.debug ({"Process file: ", path});
$display ({"Process file: ", path});
//   if (file_id == 0) log_.error ({"unable to open file ", path}); return; end
   if (file_id == 0) begin $display ({"unable to open file ", path});    return; end  //non error now ;-(
   while (! $feof (file_id)) 
     begin
	//get frst word
	string param ;
	byte c;
	string value;
	integer unused;

	unused = $fscanf (file_id, "%s", param);
	if (param.len ()) begin
`ifndef AXIOM
	   c = $fgetc (file_id);  //eat the space between symbol and value
`endif
	   unused = $fgets (value, file_id);
	   value = value.substr (0, value.len() - 2);
	end
	
//	$display ($psprintf ("got \"%s\" and \"%s\" ", param, value));

	if (param == "#include") begin
	   process_file_ (value);
	end
	else begin
	   lines_[param] = value;
//	      $display ("lines22[%s] is \"%s\"", param, lines_[param]);
	end
     end // while (! feof (file_id))
//      log_.debug ({"Completed process file: ", path});
   $display ({"Completed process file: ", path});
endtask

task dictionary_impl::read ( string path);
   process_file_ (path);
endtask


task dictionary_impl::clear ();
   lines_.delete ();
endtask

function bit dictionary_impl::put ( string name,  string value, input bit replace_existing);
  bit returned = (find (name) != "");
  if ( (! returned) || (replace_existing)) begin
    lines_[name] = value;
  end
  return returned;
endfunction

function string dictionary_impl::find ( string name); 
  string arg = teal_scan_plusargs (name);
//   $display ("%t lines \"%s\" is \"%s\" command line is \"%s\"", $time, name, lines_[name], arg);
   
  return (arg != "") ? arg : lines_[name];
endfunction

function integer dictionary_impl::find_integer ( string name, integer default_value);
   string value = find (name);
   integer returned;
   integer scan_count = 0;
   if (name != "") begin
      scan_count = $sscanf (value, "%d", returned);
   end
//   $display ("%t lines \"%s\" is \"%s\" ret is %0d", $time, name, lines_[name],  (scan_count == 1) ? returned : default_value);   
   return (scan_count == 1) ? returned : default_value;
endfunction
